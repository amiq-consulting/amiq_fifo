//----------------------------------------------------------------------
// Created by edaibr on Fri Feb 11 13:53:21 EET 2022
// Company name: amiq
// Project name: fifo
// Additional details:
// none
//----------------------------------------------------------------------

`ifndef AMIQ_FIFO_WRITE_DEFINES
`define AMIQ_FIFO_WRITE_DEFINES

// Defines for write agent
localparam M = `M;
localparam N = `N;
localparam P = `P;
`endif
